module EncoderSpeed (
    input logic CLOCK_50,
    input logic reset,
    input logic encoder_a,
    input logic encoder_b,                                                    
    output logic signed [15:0] speed
);
    // Constants
    int TIMER_MAX = 50000;

    // Internal variables for tick counting and time interval
    logic signed [15:0] tick_count, previous_tick_count;
    logic [15:0] timer;
    logic actual_A, actual_B, previous_A, previous_B;

    always_ff @(posedge CLOCK_50 or posedge reset) begin
        if (reset) begin
            tick_count <= 0;
            timer <= 0;
            speed <= 0;
            previous_A <= 0;
            previous_B <= 0;
            actual_A <= 0;
            actual_B <= 0;
        end else begin
            // Increment timer and count encoder ticks
            timer <= timer + 1;

            // Update previous states
            previous_A <= actual_A;
            previous_B <= actual_B;
            actual_A <= encoder_a;
            actual_B <= encoder_b;

            case ({previous_A, previous_B, actual_A, actual_B})
                4'b00_01, 4'b01_11, 4'b11_10, 4'b10_00: tick_count <= tick_count - 1; // Backward
                4'b00_10, 4'b10_11, 4'b11_01, 4'b01_00: tick_count <= tick_count + 1; // Forward
                default: tick_count <= tick_count;
            endcase

            // Calculate speed every TIMER_MAX cycles
            if (timer >= TIMER_MAX) begin
                speed = tick_count - previous_tick_count; // Assuming tick_count per TIMER_MAX = speed
                previous_tick_count = tick_count;
                timer <= 0;
            end
        end
    end
endmodule


module Odometer (
    input logic CLOCK_50,
    input logic reset,
    input logic encoder_a,
    input logic encoder_b,
    output logic signed [31:0] tick_count // Signed for direction
);
    logic actual_A, actual_B, previous_A, previous_B;

    always_ff @(posedge CLOCK_50 or posedge reset) begin
        if (reset) begin
            tick_count <= 0;
        end else begin
            case ({previous_A, previous_B, actual_A, actual_B})
                4'b00_01, 4'b01_11, 4'b11_10, 4'b10_00: tick_count <= tick_count - 1; // Backward
                4'b00_10, 4'b10_11, 4'b11_01, 4'b01_00: tick_count <= tick_count + 1; // Forward
                default: tick_count <= tick_count;
            endcase
            // Update previous states
            previous_A <= actual_A;
            previous_B <= actual_B;
            actual_A <= encoder_a;
            actual_B <= encoder_b;
        end
    end
endmodule




//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

module DE0_NANO_V2(

	//////////// CLOCK //////////
	input 		          		CLOCK_50,

	//////////// LED //////////
	output		     [7:0]		LED,

	//////////// KEY //////////
	input 		     [1:0]		KEY,

	//////////// EPCS //////////
	output		          		EPCS_ASDO,
	input 		          		EPCS_DATA0,
	output		          		EPCS_DCLK,
	output		          		EPCS_NCSO,

	//////////// GPIO, GPIO connect to GPIO Default //////////
	inout 		    [33:0]		GPIO,
	input 		     [1:0]		GPIO_IN
);


//========================================================
//  REG/WIRE declarations
//=======================================================


// SPI
logic 			SPI_CE, SPI_CLK, SPI_MOSI, SPI_MISO, SPI_Ready;
logic [31:0]	SPI_To_Send;
logic [7:0]		SPI_Query;
logic [3:0]		SPI_Data_Addr;
logic [31:0]	SPI_Data;
logic				SPI_Data_WE;
// Assign to external signals
assign clk = CLOCK_50;
assign reset = ~KEY[0];

assign {SPI_MOSI, SPI_CLK} = GPIO[23:22];
assign SPI_CE			   = GPIO[20];

//assign GPIO[21] = (SPI_CE) ? 1'bz : SPI_MISO;
assign GPIO[21] = SPI_MISO;
//assign SPI_To_Send = 32'hFFFFFFEC;

assign ENC_1A = GPIO[1]; // Encoder 1 Channel A
assign ENC_1B = GPIO[3]; // Encoder 1 Channel B
assign ENC_2A = GPIO[2]; // Encoder 2 Channel A
assign ENC_2B = GPIO[5]; // Encoder 2 Channel B

assign ODO_1A = GPIO[8];  // Odometer 1 Channel A
assign ODO_1B = GPIO[9];  // Odometer 1 Channel B
assign ODO_2A = GPIO[10]; // Odometer 2 Channel A
assign ODO_2B = GPIO[11]; // Odometer 2 Channel B

//=======================================================
//  Structural coding
//=======================================================
logic [7:0] address;

logic signed [15:0] left_speed, right_speed;
logic signed [31:0] left_ticks, right_ticks;


// SPI slave
spi_slave spi(
	.SPI_CLK(SPI_CLK),
	.SPI_CS(SPI_CE),
	.SPI_MOSI(SPI_MOSI),
	.clk(clk),
	.SPI_MISO(SPI_MISO),
	.ToSend(SPI_To_Send),
	.Query(SPI_Query),
	.Ready(SPI_Ready),
	.DataAddr(SPI_Data_Addr),
	.Data(SPI_Data),
	.Data_WE(SPI_Data_WE),
    );


 // Instantiate modules
    EncoderSpeed left_encoder_speed (
        .CLOCK_50(clk), .reset(reset), 
        .encoder_a(ENC_1A), .encoder_b(ENC_1B), 
        .speed(left_speed)
    );

    EncoderSpeed right_encoder_speed (
        .CLOCK_50(clk), .reset(reset), 
        .encoder_a(ENC_2A), .encoder_b(ENC_2B), 
        .speed(right_speed)
    );

    Odometer left_odometer (
        .CLOCK_50(clk), .reset(reset), 
        .encoder_a(ODO_1A), .encoder_b(ODO_1B), 
        .tick_count(left_ticks)
    );

    Odometer right_odometer (
        .CLOCK_50(clk), .reset(reset), 
        .encoder_a(ODO_2A), .encoder_b(ODO_2B), 
        .tick_count(right_ticks)
    );

assign SPI_To_Send = left_speed;

/*always  begin

		address <= SPI_Query;
		
		case (address)
			8'h10: SPI_To_Send = left_speed;
			8'h11: SPI_To_Send = right_speed;
			8'h12: SPI_To_Send = left_ticks;
			8'h13: SPI_To_Send = right_ticks;
			// 8'h7F in decimal is 127
			8'h7F: SPI_To_Send = 32'd127;
		endcase
	end
*/

assign LED = SPI_To_Send[7:0];

endmodule
