module EncoderSpeed (
    input logic CLOCK_50,
    input logic reset,
    input logic encoder_a,
    input logic encoder_b,                                                    
    output logic signed [31:0] speed
);
    // Constants
    int TIMER_MAX = 500000;

    // Internal variables for tick counting and time interval
    logic signed [31:0] tick_count;
    logic [31:0] timer;
    logic actual_A, actual_B, previous_A, previous_B;

    always_ff @(posedge CLOCK_50 or posedge reset) begin
        if (reset) begin
            tick_count <= 0;
            timer <= 0;
            speed <= 0;
        end else begin
            // Increment timer and count encoder ticks
            timer <= timer + 1;

            // Update previous states
            previous_A <= actual_A;
            previous_B <= actual_B;
            actual_A <= encoder_a;
            actual_B <= encoder_b;

            case ({previous_A, previous_B, actual_A, actual_B})
                4'b00_01, 4'b01_11, 4'b11_10, 4'b10_00: tick_count <= tick_count + 1; // Forward
                4'b00_10, 4'b10_11, 4'b11_01, 4'b01_00: tick_count <= tick_count - 1; // Backward
                default: tick_count <= tick_count;
            endcase

            // Calculate speed every TIMER_MAX cycles
            if (timer >= TIMER_MAX) begin
                speed <= tick_count; // Assuming tick_count per TIMER_MAX = speed
                tick_count <= 0;
                timer <= 0;
            end

            

        end
    end
endmodule


module Odometer (
    input logic CLOCK_50,
    input logic reset,
    input logic encoder_a,
    input logic encoder_b,
    output logic signed [31:0] tick_count // Signed for direction
);
    logic actual_A, actual_B, previous_A, previous_B;

    always_ff @(posedge CLOCK_50 or posedge reset) begin
        if (reset) begin
            tick_count <= 0;
        end else begin
            case ({previous_A, previous_B, actual_A, actual_B})
                4'b00_01, 4'b01_11, 4'b11_10, 4'b10_00: tick_count <= tick_count - 1; // Backward
                4'b00_10, 4'b10_11, 4'b11_01, 4'b01_00: tick_count <= tick_count + 1; // Forward
                default: tick_count <= tick_count;
            endcase
            // Update previous states
            previous_A <= actual_A;
            previous_B <= actual_B;
            actual_A <= encoder_a;
            actual_B <= encoder_b;
        end
    end
endmodule




//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

module DE0_NANO_V3(

	//////////// CLOCK //////////
	input 		          		CLOCK_50,

	//////////// LED //////////
	output		     [7:0]		LED,

	//////////// KEY //////////
	input 		     [1:0]		KEY,

	//////////// SW //////////
	input 		     [3:0]		SW,

	//////////// SDRAM //////////
	output		    [12:0]		DRAM_ADDR,
	output		     [1:0]		DRAM_BA,
	output		          		DRAM_CAS_N,
	output		          		DRAM_CKE,
	output		          		DRAM_CLK,
	output		          		DRAM_CS_N,
	inout 		    [15:0]		DRAM_DQ,
	output		     [1:0]		DRAM_DQM,
	output		          		DRAM_RAS_N,
	output		          		DRAM_WE_N,

	//////////// EPCS //////////
	output		          		EPCS_ASDO,
	input 		          		EPCS_DATA0,
	output		          		EPCS_DCLK,
	output		          		EPCS_NCSO,

	//////////// Accelerometer and EEPROM //////////
	output		          		G_SENSOR_CS_N,
	input 		          		G_SENSOR_INT,
	output		          		I2C_SCLK,
	inout 		          		I2C_SDAT,

	//////////// ADC //////////
	output		          		ADC_CS_N,
	output		          		ADC_SADDR,
	output		          		ADC_SCLK,
	input 		          		ADC_SDAT,

	//////////// GPIO_0, GPIO_0 connect to GPIO Default //////////
	inout 		    [33:0]		GPIO_1,
	input 		     [1:0]		GPIO_1_IN,

	//////////// GPIO_1, GPIO_1 connect to GPIO Default //////////
	inout 		    [33:0]		GPIO_2,
	input 		     [1:0]		GPIO_2_IN
);


//=======================================================
//  REG/WIRE declarations
//=======================================================

// SPI
logic 			SPI_CE, SPI_CLK, SPI_MOSI, SPI_MISO, SPI_Ready;
logic [31:0]	SPI_To_Send;
logic [7:0]		SPI_Query;
logic [3:0]		SPI_Data_Addr;
logic [31:0]	SPI_Data;
logic				SPI_Data_WE;
// Assign to external signals
assign clk = CLOCK_50;
logic internal_reset;
assign reset = ~KEY[0] | internal_reset;

assign SPI_MOSI = GPIO_2_IN[1];
assign SPI_MISO = (SPI_CE) ? 1'bz : GPIO_2[1];
assign SPI_CLK  = GPIO_2[2];
assign SPI_CE   = GPIO_2[4];
//assign SPI_To_Send = 32'hFFFFFFEC; to debug SPI if needed

assign ENC_1A = GPIO_2[10]; // Encoder 1 Channel A
assign ENC_1B = GPIO_2[12]; // Encoder 1 Channel B
assign ENC_2A = GPIO_2[16]; // Encoder 2 Channel A
assign ENC_2B = GPIO_2[18]; // Encoder 2 Channel B

assign ODO_1A = GPIO_2[22];  // Odometer 1 Channel A
assign ODO_1B = GPIO_2[24];  // Odometer 1 Channel B
assign ODO_2A = GPIO_2[28]; // Odometer 2 Channel A
assign ODO_2B = GPIO_2[30]; // Odometer 2 Channel B

//=======================================================
//  Structural coding
//=======================================================
logic [7:0] address;

logic signed [31:0] left_speed, right_speed;
logic signed [31:0] left_ticks, right_ticks;


// SPI slave
spi_slave spi(
	.SPI_CLK(SPI_CLK),
	.SPI_CS(SPI_CE),
	.SPI_MOSI(SPI_MOSI),
	.clk(clk),
	.SPI_MISO(SPI_MISO),
	.ToSend(SPI_To_Send),
	.Query(SPI_Query),
	.Ready(SPI_Ready),
	.DataAddr(SPI_Data_Addr),
	.Data(SPI_Data),
	.Data_WE(SPI_Data_WE),
    );


 // Instantiate modules
    EncoderSpeed left_encoder_speed (
        .CLOCK_50(clk), .reset(reset), 
        .encoder_a(ENC_1A), .encoder_b(ENC_1B), 
        .speed(left_speed)
    );

    EncoderSpeed right_encoder_speed (
        .CLOCK_50(clk), .reset(reset), 
        .encoder_a(ENC_2A), .encoder_b(ENC_2B), 
        .speed(right_speed)
    );

    Odometer left_odometer (
        .CLOCK_50(clk), .reset(reset), 
        .encoder_a(ODO_1A), .encoder_b(ODO_1B), 
        .tick_count(left_ticks)
    );

    Odometer right_odometer (
        .CLOCK_50(clk), .reset(reset), 
        .encoder_a(ODO_2A), .encoder_b(ODO_2B), 
        .tick_count(right_ticks)
    );

always_ff @(posedge SPI_Ready) begin
    //address = SPI_Query;
    case (SPI_Query)
        8'h10: SPI_To_Send <= left_speed;
        8'h11: SPI_To_Send <= -right_speed;
        8'h12: SPI_To_Send <= -left_ticks;
        8'h13: SPI_To_Send <= right_ticks;
        8'h7F: ; // Do nothing for reset query
        default: SPI_To_Send <= SPI_To_Send; // Hold previous value
    endcase
end


// Generate a one-clock-cycle pulse for `internal_reset`
always_ff @(posedge clk) begin
    if (SPI_Query == 8'h7F) begin
        internal_reset <= 1;
    end else begin
        internal_reset <= 0;
    end
end



assign LED = right_ticks[7:0];

endmodule
